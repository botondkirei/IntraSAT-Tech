-- utils package to be used in wisat2 project
-- Company : UTCN
-- Employee : Kirei Botond
-- Rev - 0.01 -file created

library IEEE;
use IEEE.std_logic_1164.all;

package utils is
	type SpWIO is record
	end record;
	type FMCIO is record
	end record;
end package;

package body utils is
end package body;
